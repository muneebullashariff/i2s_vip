// basic file added
